library ieee;
use ieee.std_logic_1164.all;

entity dpram is
    generic
    (
        mem_size    : natural := 95 * 95;
        data_width  : natural := 8
    );
   port 
   (   
        i_clk_a        : in std_logic;
        i_clk_b        : in std_logic;

        i_data_a    : in std_logic_vector(data_width-1 downto 0);
        i_data_b    : in std_logic_vector(data_width-1 downto 0);
        i_addr_a    : in natural range 0 to mem_size-1;
        i_addr_b    : in natural range 0 to mem_size-1;
        i_we_a      : in std_logic := '1';
        i_we_b      : in std_logic := '1';
        o_q_a       : out std_logic_vector(data_width-1 downto 0);
        o_q_b       : out std_logic_vector(data_width-1 downto 0)
   );
   
end dpram;

architecture rtl of dpram is
    -- Build a 2-D array type for the RAM
    subtype word_t is std_logic_vector(data_width-1 downto 0);
    type memory_t is array(0 to mem_size-1) of word_t;
    
    -- Declare the RAM
    shared variable ram : memory_t := (
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"da", x"ff", x"ff", x"ff", 
        x"b5", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"53", 
        x"ff", x"ff", x"ff", x"84", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"6c", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"b5", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"9d", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"ff", x"ff", x"ff", x"53", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ce", x"ff", x"da", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"ff", x"53", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ce", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"f3", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"f3", x"ff", x"ff", 
        x"ff", x"ff", x"78", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"90", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"da", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"78", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ce", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"b5", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"f3", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"90", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"90", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"3a", x"3a", x"5f", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"3a", x"46", x"46", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"3a", 
        x"6c", x"c2", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"46", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"3a", x"a9", x"ff", x"f3", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"6c", x"ff", x"ff", x"ff", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"f3", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"78", x"ff", x"ff", x"ff", x"3a", x"ff", x"ff", x"ff", x"ff", x"c2", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"6c", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"78", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"ff", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ce", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"3a", x"3a", x"9d", x"6c", x"3a", x"3a", x"3a", x"3a", x"9d", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"f3", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"84", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"84", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"c2", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"84", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ce", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"ff", x"ce", x"6c", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"9d", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"78", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"c2", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"5f", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"da", x"3a", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"e6", 
        x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", x"ff", x"ff", x"ff", 
        x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ce", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"84", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"53", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", 
        x"ff", x"3a", x"84", x"ff", x"ff", x"ff", x"90", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ce", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ce", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"f3", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"da", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"46", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"46", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"b5", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"ff", x"ff", x"ff", x"ff", x"46", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", 
        x"3a", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"6c", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
        x"ff", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff", x"3a", x"3a", 
        x"3a", x"3a", x"3a", x"3a", x"3a", x"3a", x"ff", x"ff", x"ff", x"ff"
    );
begin
    -- Port A
    process(i_clk_a)
    begin
        if(rising_edge(i_clk_a)) then 
            if(i_we_a = '1') then
                ram(i_addr_a) := i_data_a;
            end if;
            o_q_a <= ram(i_addr_a);
        end if;
    end process;
    
    -- Port B
    process(i_clk_b)
    begin
        if(rising_edge(i_clk_b)) then
            if(i_we_b = '1') then
                ram(i_addr_b) := i_data_b;
            end if;
            o_q_b <= ram(i_addr_b);
        end if;
    end process;
end rtl;
